module template
(
        input wire clk,
        input wire rst
);

always @(posedge clk)
begin
        if (rst)
        begin

        end else
        begin

        end
end

endmodule
